// Copyright 2016 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


interface vgm_wb_master_interface(input bit RST_I, input bit CLK_I);
  logic CYC_O;
  logic STB_O;
  logic WE_O;
  logic [31:0] ADR_O;
  logic [31:0] DAT_O;

  logic ACK_I;
  logic [31:0] DAT_I;
endinterface
